module redis

// https://github.com/vlang/v/issues/18900
// Once this bug is fixed, replace json2.Any with this type
interface Any {}
