module redis

interface Any {}
